/*ģ��˵��
ʱ�ӣ�50M�ķ�Ƶ����12.5M

*/
module dac_c (
    //global clock
    input  clk,
    input  rst_n,

    //user interface
    output sclk

);
//adc��ʱ��
//---------------------------------------------------------------------
    //������
    always @(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            cnt <= 0;
          end
        else if(add_cnt)begin
          if(end_cnt)
             cnt <= 0;
          else
             cnt <= cnt + 1;
          end      
    end

    assign add_cnt = ;
    assign end_cnt = add_cnt && cnt == ;

    //����adc
    always  @(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            sclk <= 1;
        end
        else if(end_cnt)begin
            sclk <= !sclk;
        end
    end
//---------------------------------------------------------------------



endmodule